module image(input [4:0] x, input [4:0] y, output reg [7:0] r, output reg [7:0] g, output reg [7:0] b);
wire [9:0] ix = x << 5 | y;
always @(ix) begin
case(ix)
	10'h000: begin r = 8'h90; g = 8'hac; b = 8'haa; end
	10'h020: begin r = 8'h94; g = 8'hac; b = 8'haa; end
	10'h040: begin r = 8'h93; g = 8'haa; b = 8'ha7; end
	10'h060: begin r = 8'h95; g = 8'hab; b = 8'haa; end
	10'h080: begin r = 8'h95; g = 8'hab; b = 8'ha9; end
	10'h0a0: begin r = 8'h94; g = 8'hab; b = 8'ha9; end
	10'h0c0: begin r = 8'h95; g = 8'had; b = 8'haa; end
	10'h0e0: begin r = 8'h96; g = 8'hac; b = 8'hae; end
	10'h100: begin r = 8'h98; g = 8'had; b = 8'hae; end
	10'h120: begin r = 8'h97; g = 8'hac; b = 8'had; end
	10'h140: begin r = 8'h94; g = 8'haa; b = 8'hac; end
	10'h160: begin r = 8'h93; g = 8'ha9; b = 8'had; end
	10'h180: begin r = 8'h90; g = 8'ha8; b = 8'ha9; end
	10'h1a0: begin r = 8'h98; g = 8'hac; b = 8'ha7; end
	10'h1c0: begin r = 8'hb1; g = 8'hba; b = 8'hb2; end
	10'h1e0: begin r = 8'hc8; g = 8'hca; b = 8'hbc; end
	10'h200: begin r = 8'hd5; g = 8'hd3; b = 8'hc7; end
	10'h220: begin r = 8'hd6; g = 8'hd8; b = 8'hc6; end
	10'h240: begin r = 8'hcc; g = 8'hce; b = 8'hc1; end
	10'h260: begin r = 8'hb2; g = 8'hbf; b = 8'hb6; end
	10'h280: begin r = 8'h95; g = 8'ha7; b = 8'h9f; end
	10'h2a0: begin r = 8'h87; g = 8'h9d; b = 8'h99; end
	10'h2c0: begin r = 8'h89; g = 8'h9d; b = 8'h9c; end
	10'h2e0: begin r = 8'h89; g = 8'h9d; b = 8'h9e; end
	10'h300: begin r = 8'h86; g = 8'h9c; b = 8'h9d; end
	10'h320: begin r = 8'h85; g = 8'h9b; b = 8'h99; end
	10'h340: begin r = 8'h82; g = 8'h98; b = 8'h94; end
	10'h360: begin r = 8'h82; g = 8'h99; b = 8'h91; end
	10'h380: begin r = 8'h80; g = 8'h95; b = 8'h91; end
	10'h3a0: begin r = 8'h80; g = 8'h95; b = 8'h94; end
	10'h3c0: begin r = 8'h8a; g = 8'h9c; b = 8'h9e; end
	10'h3e0: begin r = 8'h85; g = 8'h94; b = 8'h97; end
	10'h001: begin r = 8'h90; g = 8'hae; b = 8'had; end
	10'h021: begin r = 8'h93; g = 8'had; b = 8'hab; end
	10'h041: begin r = 8'h95; g = 8'had; b = 8'haa; end
	10'h061: begin r = 8'h97; g = 8'had; b = 8'hac; end
	10'h081: begin r = 8'h96; g = 8'hac; b = 8'had; end
	10'h0a1: begin r = 8'h98; g = 8'had; b = 8'hae; end
	10'h0c1: begin r = 8'h98; g = 8'hae; b = 8'hae; end
	10'h0e1: begin r = 8'h98; g = 8'had; b = 8'hae; end
	10'h101: begin r = 8'h9a; g = 8'hb0; b = 8'hb1; end
	10'h121: begin r = 8'h99; g = 8'hae; b = 8'haf; end
	10'h141: begin r = 8'h94; g = 8'hab; b = 8'hac; end
	10'h161: begin r = 8'h9d; g = 8'hb1; b = 8'hac; end
	10'h181: begin r = 8'hbd; g = 8'hc0; b = 8'hb7; end
	10'h1a1: begin r = 8'hc7; g = 8'hc2; b = 8'hb2; end
	10'h1c1: begin r = 8'hc7; g = 8'hbd; b = 8'ha8; end
	10'h1e1: begin r = 8'hc1; g = 8'hb5; b = 8'h9b; end
	10'h201: begin r = 8'hc9; g = 8'hbb; b = 8'ha5; end
	10'h221: begin r = 8'hcf; g = 8'hc0; b = 8'ha8; end
	10'h241: begin r = 8'hd4; g = 8'hc2; b = 8'ha6; end
	10'h261: begin r = 8'hd7; g = 8'hcd; b = 8'hb1; end
	10'h281: begin r = 8'he2; g = 8'hdf; b = 8'hcb; end
	10'h2a1: begin r = 8'hd0; g = 8'hd5; b = 8'hc8; end
	10'h2c1: begin r = 8'h94; g = 8'ha6; b = 8'ha0; end
	10'h2e1: begin r = 8'h8b; g = 8'ha1; b = 8'h9f; end
	10'h301: begin r = 8'h8a; g = 8'h9f; b = 8'h9f; end
	10'h321: begin r = 8'h89; g = 8'h9e; b = 8'h9f; end
	10'h341: begin r = 8'h86; g = 8'h9d; b = 8'h99; end
	10'h361: begin r = 8'h84; g = 8'h9b; b = 8'h97; end
	10'h381: begin r = 8'h83; g = 8'h98; b = 8'h97; end
	10'h3a1: begin r = 8'h82; g = 8'h97; b = 8'h97; end
	10'h3c1: begin r = 8'h7f; g = 8'h93; b = 8'h94; end
	10'h3e1: begin r = 8'h82; g = 8'h94; b = 8'h96; end
	10'h002: begin r = 8'h91; g = 8'hae; b = 8'hae; end
	10'h022: begin r = 8'h96; g = 8'hb0; b = 8'haf; end
	10'h042: begin r = 8'h97; g = 8'hb0; b = 8'hb0; end
	10'h062: begin r = 8'h97; g = 8'haf; b = 8'haf; end
	10'h082: begin r = 8'h96; g = 8'had; b = 8'had; end
	10'h0a2: begin r = 8'h98; g = 8'had; b = 8'hae; end
	10'h0c2: begin r = 8'h99; g = 8'hae; b = 8'haf; end
	10'h0e2: begin r = 8'h98; g = 8'hae; b = 8'haf; end
	10'h102: begin r = 8'h97; g = 8'haf; b = 8'hb1; end
	10'h122: begin r = 8'h9a; g = 8'hb0; b = 8'haf; end
	10'h142: begin r = 8'hb4; g = 8'hbd; b = 8'hb4; end
	10'h162: begin r = 8'hae; g = 8'ha8; b = 8'h92; end
	10'h182: begin r = 8'h7f; g = 8'h6e; b = 8'h4b; end
	10'h1a2: begin r = 8'h6d; g = 8'h59; b = 8'h36; end
	10'h1c2: begin r = 8'h74; g = 8'h5f; b = 8'h43; end
	10'h1e2: begin r = 8'h87; g = 8'h73; b = 8'h55; end
	10'h202: begin r = 8'h97; g = 8'h86; b = 8'h67; end
	10'h222: begin r = 8'h9a; g = 8'h88; b = 8'h6a; end
	10'h242: begin r = 8'ha6; g = 8'h95; b = 8'h73; end
	10'h262: begin r = 8'hb5; g = 8'ha3; b = 8'h7f; end
	10'h282: begin r = 8'hb9; g = 8'ha4; b = 8'h84; end
	10'h2a2: begin r = 8'hc2; g = 8'hb3; b = 8'h9b; end
	10'h2c2: begin r = 8'he7; g = 8'he3; b = 8'hd1; end
	10'h2e2: begin r = 8'hab; g = 8'hb9; b = 8'hac; end
	10'h302: begin r = 8'h90; g = 8'ha3; b = 8'ha1; end
	10'h322: begin r = 8'h8c; g = 8'ha2; b = 8'ha0; end
	10'h342: begin r = 8'h89; g = 8'h9f; b = 8'h9e; end
	10'h362: begin r = 8'h85; g = 8'h9b; b = 8'h99; end
	10'h382: begin r = 8'h87; g = 8'h9b; b = 8'h9c; end
	10'h3a2: begin r = 8'h86; g = 8'h9c; b = 8'h9d; end
	10'h3c2: begin r = 8'h83; g = 8'h97; b = 8'h98; end
	10'h3e2: begin r = 8'h84; g = 8'h96; b = 8'h96; end
	10'h003: begin r = 8'h91; g = 8'haf; b = 8'hb1; end
	10'h023: begin r = 8'h95; g = 8'hb2; b = 8'hb5; end
	10'h043: begin r = 8'h97; g = 8'hb0; b = 8'hb3; end
	10'h063: begin r = 8'h97; g = 8'haf; b = 8'hb2; end
	10'h083: begin r = 8'h98; g = 8'hb0; b = 8'hb0; end
	10'h0a3: begin r = 8'h97; g = 8'hb0; b = 8'hb0; end
	10'h0c3: begin r = 8'h97; g = 8'haf; b = 8'haf; end
	10'h0e3: begin r = 8'h96; g = 8'hb0; b = 8'haf; end
	10'h103: begin r = 8'h98; g = 8'hb2; b = 8'hb0; end
	10'h123: begin r = 8'h9b; g = 8'h97; b = 8'h87; end
	10'h143: begin r = 8'h94; g = 8'h7b; b = 8'h55; end
	10'h163: begin r = 8'hac; g = 8'h87; b = 8'h4c; end
	10'h183: begin r = 8'hbb; g = 8'h8b; b = 8'h3e; end
	10'h1a3: begin r = 8'hb7; g = 8'h8a; b = 8'h46; end
	10'h1c3: begin r = 8'hab; g = 8'h85; b = 8'h51; end
	10'h1e3: begin r = 8'h9b; g = 8'h84; b = 8'h5c; end
	10'h203: begin r = 8'ha8; g = 8'h8b; b = 8'h62; end
	10'h223: begin r = 8'hb6; g = 8'ha1; b = 8'h83; end
	10'h243: begin r = 8'hbd; g = 8'ha8; b = 8'h87; end
	10'h263: begin r = 8'hc4; g = 8'hac; b = 8'h8d; end
	10'h283: begin r = 8'hce; g = 8'hb5; b = 8'h97; end
	10'h2a3: begin r = 8'hdb; g = 8'hc5; b = 8'had; end
	10'h2c3: begin r = 8'hc7; g = 8'hb4; b = 8'h9e; end
	10'h2e3: begin r = 8'hdc; g = 8'hd1; b = 8'hbe; end
	10'h303: begin r = 8'hb5; g = 8'hbf; b = 8'hb9; end
	10'h323: begin r = 8'h8f; g = 8'ha5; b = 8'ha3; end
	10'h343: begin r = 8'h8a; g = 8'ha2; b = 8'ha3; end
	10'h363: begin r = 8'h87; g = 8'ha0; b = 8'h9d; end
	10'h383: begin r = 8'h8b; g = 8'ha0; b = 8'ha1; end
	10'h3a3: begin r = 8'h88; g = 8'h9d; b = 8'h9e; end
	10'h3c3: begin r = 8'h88; g = 8'h9d; b = 8'h9e; end
	10'h3e3: begin r = 8'h86; g = 8'h9b; b = 8'h9a; end
	10'h004: begin r = 8'h93; g = 8'hb1; b = 8'hb3; end
	10'h024: begin r = 8'h94; g = 8'hb2; b = 8'hb4; end
	10'h044: begin r = 8'h96; g = 8'hb1; b = 8'hb4; end
	10'h064: begin r = 8'h98; g = 8'hb0; b = 8'hb4; end
	10'h084: begin r = 8'h97; g = 8'haf; b = 8'hb2; end
	10'h0a4: begin r = 8'h97; g = 8'hb0; b = 8'hb2; end
	10'h0c4: begin r = 8'h95; g = 8'had; b = 8'had; end
	10'h0e4: begin r = 8'h94; g = 8'hac; b = 8'hac; end
	10'h104: begin r = 8'h71; g = 8'h6e; b = 8'h64; end
	10'h124: begin r = 8'h7b; g = 8'h61; b = 8'h38; end
	10'h144: begin r = 8'hb6; g = 8'h8c; b = 8'h45; end
	10'h164: begin r = 8'hca; g = 8'h99; b = 8'h45; end
	10'h184: begin r = 8'hd3; g = 8'h9e; b = 8'h45; end
	10'h1a4: begin r = 8'hd8; g = 8'ha2; b = 8'h56; end
	10'h1c4: begin r = 8'hd9; g = 8'ha6; b = 8'h55; end
	10'h1e4: begin r = 8'hd9; g = 8'haa; b = 8'h61; end
	10'h204: begin r = 8'hcd; g = 8'ha7; b = 8'h6d; end
	10'h224: begin r = 8'hd0; g = 8'hae; b = 8'h7d; end
	10'h244: begin r = 8'hdc; g = 8'hba; b = 8'h99; end
	10'h264: begin r = 8'he0; g = 8'hbe; b = 8'h9f; end
	10'h284: begin r = 8'he6; g = 8'hc4; b = 8'ha9; end
	10'h2a4: begin r = 8'he1; g = 8'hbf; b = 8'h9c; end
	10'h2c4: begin r = 8'hd7; g = 8'hb1; b = 8'h8b; end
	10'h2e4: begin r = 8'hcf; g = 8'hb1; b = 8'h8e; end
	10'h304: begin r = 8'hd1; g = 8'hc6; b = 8'hb5; end
	10'h324: begin r = 8'h98; g = 8'ha8; b = 8'ha4; end
	10'h344: begin r = 8'h8a; g = 8'ha3; b = 8'ha0; end
	10'h364: begin r = 8'h89; g = 8'ha1; b = 8'ha1; end
	10'h384: begin r = 8'h8a; g = 8'h9e; b = 8'h9f; end
	10'h3a4: begin r = 8'h87; g = 8'h9e; b = 8'h9e; end
	10'h3c4: begin r = 8'h86; g = 8'h9b; b = 8'h9c; end
	10'h3e4: begin r = 8'h86; g = 8'h9a; b = 8'h9b; end
	10'h005: begin r = 8'h94; g = 8'hb1; b = 8'hb4; end
	10'h025: begin r = 8'h96; g = 8'hb4; b = 8'hb6; end
	10'h045: begin r = 8'h97; g = 8'hb5; b = 8'hb7; end
	10'h065: begin r = 8'h99; g = 8'hb1; b = 8'hb5; end
	10'h085: begin r = 8'h98; g = 8'hb0; b = 8'hb0; end
	10'h0a5: begin r = 8'h98; g = 8'haf; b = 8'haf; end
	10'h0c5: begin r = 8'h94; g = 8'hac; b = 8'hab; end
	10'h0e5: begin r = 8'h75; g = 8'h79; b = 8'h69; end
	10'h105: begin r = 8'h83; g = 8'h71; b = 8'h55; end
	10'h125: begin r = 8'haf; g = 8'h87; b = 8'h4b; end
	10'h145: begin r = 8'hd3; g = 8'h9a; b = 8'h4b; end
	10'h165: begin r = 8'hd5; g = 8'ha0; b = 8'h47; end
	10'h185: begin r = 8'hde; g = 8'ha6; b = 8'h55; end
	10'h1a5: begin r = 8'he5; g = 8'hab; b = 8'h62; end
	10'h1c5: begin r = 8'he9; g = 8'hb0; b = 8'h68; end
	10'h1e5: begin r = 8'he9; g = 8'haf; b = 8'h66; end
	10'h205: begin r = 8'he9; g = 8'hb0; b = 8'h6b; end
	10'h225: begin r = 8'he2; g = 8'hb0; b = 8'h6f; end
	10'h245: begin r = 8'hdf; g = 8'haf; b = 8'h79; end
	10'h265: begin r = 8'he0; g = 8'hb4; b = 8'h84; end
	10'h285: begin r = 8'he8; g = 8'hba; b = 8'h95; end
	10'h2a5: begin r = 8'he3; g = 8'hb5; b = 8'h84; end
	10'h2c5: begin r = 8'hd5; g = 8'hab; b = 8'h6d; end
	10'h2e5: begin r = 8'hce; g = 8'ha6; b = 8'h69; end
	10'h305: begin r = 8'hcd; g = 8'hb1; b = 8'h8c; end
	10'h325: begin r = 8'hb0; g = 8'hae; b = 8'h9f; end
	10'h345: begin r = 8'h8e; g = 8'ha1; b = 8'h9a; end
	10'h365: begin r = 8'h88; g = 8'ha1; b = 8'h9d; end
	10'h385: begin r = 8'h85; g = 8'h9e; b = 8'h9e; end
	10'h3a5: begin r = 8'h84; g = 8'h9c; b = 8'h9d; end
	10'h3c5: begin r = 8'h86; g = 8'h9b; b = 8'h9c; end
	10'h3e5: begin r = 8'h83; g = 8'h9b; b = 8'h9b; end
	10'h006: begin r = 8'h95; g = 8'hb3; b = 8'hb5; end
	10'h026: begin r = 8'h97; g = 8'hb5; b = 8'hb7; end
	10'h046: begin r = 8'h98; g = 8'hb4; b = 8'hb7; end
	10'h066: begin r = 8'h9a; g = 8'hb2; b = 8'hb7; end
	10'h086: begin r = 8'h99; g = 8'hb0; b = 8'hb1; end
	10'h0a6: begin r = 8'h98; g = 8'hae; b = 8'had; end
	10'h0c6: begin r = 8'h8b; g = 8'h98; b = 8'h92; end
	10'h0e6: begin r = 8'ha0; g = 8'h97; b = 8'h83; end
	10'h106: begin r = 8'ha4; g = 8'h8d; b = 8'h69; end
	10'h126: begin r = 8'hc7; g = 8'h98; b = 8'h48; end
	10'h146: begin r = 8'hd5; g = 8'h9e; b = 8'h4e; end
	10'h166: begin r = 8'hd7; g = 8'ha0; b = 8'h4f; end
	10'h186: begin r = 8'he2; g = 8'ha9; b = 8'h62; end
	10'h1a6: begin r = 8'he9; g = 8'had; b = 8'h70; end
	10'h1c6: begin r = 8'hf4; g = 8'hb8; b = 8'h81; end
	10'h1e6: begin r = 8'hf7; g = 8'hbc; b = 8'h86; end
	10'h206: begin r = 8'hf4; g = 8'hba; b = 8'h80; end
	10'h226: begin r = 8'hf3; g = 8'hb7; b = 8'h7d; end
	10'h246: begin r = 8'hf3; g = 8'hbb; b = 8'h81; end
	10'h266: begin r = 8'hf3; g = 8'hb9; b = 8'h80; end
	10'h286: begin r = 8'hf9; g = 8'hbf; b = 8'h8b; end
	10'h2a6: begin r = 8'hf1; g = 8'hbc; b = 8'h85; end
	10'h2c6: begin r = 8'hea; g = 8'hb6; b = 8'h7f; end
	10'h2e6: begin r = 8'hdc; g = 8'hb2; b = 8'h7d; end
	10'h306: begin r = 8'hd1; g = 8'ha9; b = 8'h78; end
	10'h326: begin r = 8'hc4; g = 8'haa; b = 8'h8b; end
	10'h346: begin r = 8'haf; g = 8'had; b = 8'ha1; end
	10'h366: begin r = 8'h8a; g = 8'ha4; b = 8'h9d; end
	10'h386: begin r = 8'h85; g = 8'ha3; b = 8'h9f; end
	10'h3a6: begin r = 8'h86; g = 8'ha1; b = 8'ha0; end
	10'h3c6: begin r = 8'h87; g = 8'h9f; b = 8'h9f; end
	10'h3e6: begin r = 8'h85; g = 8'h9d; b = 8'h9d; end
	10'h007: begin r = 8'h99; g = 8'hb4; b = 8'hb7; end
	10'h027: begin r = 8'h97; g = 8'hb5; b = 8'hb7; end
	10'h047: begin r = 8'h99; g = 8'hb4; b = 8'hb7; end
	10'h067: begin r = 8'h9c; g = 8'hb3; b = 8'hb7; end
	10'h087: begin r = 8'h9a; g = 8'hb2; b = 8'hb2; end
	10'h0a7: begin r = 8'h95; g = 8'hac; b = 8'haa; end
	10'h0c7: begin r = 8'h6e; g = 8'h6c; b = 8'h5d; end
	10'h0e7: begin r = 8'h94; g = 8'h86; b = 8'h6c; end
	10'h107: begin r = 8'ha9; g = 8'h85; b = 8'h43; end
	10'h127: begin r = 8'hd6; g = 8'ha2; b = 8'h49; end
	10'h147: begin r = 8'hd5; g = 8'ha1; b = 8'h4e; end
	10'h167: begin r = 8'hda; g = 8'ha2; b = 8'h56; end
	10'h187: begin r = 8'he0; g = 8'ha8; b = 8'h5e; end
	10'h1a7: begin r = 8'heb; g = 8'hb1; b = 8'h71; end
	10'h1c7: begin r = 8'hfc; g = 8'hc1; b = 8'h8c; end
	10'h1e7: begin r = 8'hfd; g = 8'hcf; b = 8'ha4; end
	10'h207: begin r = 8'hfe; g = 8'hc7; b = 8'h98; end
	10'h227: begin r = 8'hf9; g = 8'hbb; b = 8'h84; end
	10'h247: begin r = 8'hf6; g = 8'hb8; b = 8'h7f; end
	10'h267: begin r = 8'hfc; g = 8'hbb; b = 8'h85; end
	10'h287: begin r = 8'hff; g = 8'hc5; b = 8'h95; end
	10'h2a7: begin r = 8'hfe; g = 8'hc3; b = 8'h93; end
	10'h2c7: begin r = 8'hf7; g = 8'hc0; b = 8'h96; end
	10'h2e7: begin r = 8'hf3; g = 8'hc1; b = 8'h97; end
	10'h307: begin r = 8'hdd; g = 8'hb0; b = 8'h81; end
	10'h327: begin r = 8'hd1; g = 8'ha9; b = 8'h7c; end
	10'h347: begin r = 8'hbb; g = 8'ha8; b = 8'h91; end
	10'h367: begin r = 8'ha3; g = 8'hb0; b = 8'ha8; end
	10'h387: begin r = 8'h87; g = 8'ha5; b = 8'ha4; end
	10'h3a7: begin r = 8'h8c; g = 8'ha7; b = 8'ha6; end
	10'h3c7: begin r = 8'h8c; g = 8'ha4; b = 8'ha4; end
	10'h3e7: begin r = 8'h89; g = 8'ha1; b = 8'ha1; end
	10'h008: begin r = 8'h9a; g = 8'hb5; b = 8'hb8; end
	10'h028: begin r = 8'h9b; g = 8'hb3; b = 8'hb7; end
	10'h048: begin r = 8'h9b; g = 8'hb3; b = 8'hb7; end
	10'h068: begin r = 8'h9a; g = 8'hb3; b = 8'hb7; end
	10'h088: begin r = 8'h96; g = 8'hb2; b = 8'hb4; end
	10'h0a8: begin r = 8'h8f; g = 8'ha0; b = 8'h9e; end
	10'h0c8: begin r = 8'h86; g = 8'h7c; b = 8'h6d; end
	10'h0e8: begin r = 8'h96; g = 8'h81; b = 8'h68; end
	10'h108: begin r = 8'hc3; g = 8'h8d; b = 8'h44; end
	10'h128: begin r = 8'hd5; g = 8'ha3; b = 8'h4f; end
	10'h148: begin r = 8'hd1; g = 8'h9d; b = 8'h47; end
	10'h168: begin r = 8'hdb; g = 8'ha3; b = 8'h56; end
	10'h188: begin r = 8'hdf; g = 8'ha5; b = 8'h57; end
	10'h1a8: begin r = 8'he7; g = 8'hae; b = 8'h6a; end
	10'h1c8: begin r = 8'hf0; g = 8'hbb; b = 8'h86; end
	10'h1e8: begin r = 8'hfd; g = 8'hcf; b = 8'ha6; end
	10'h208: begin r = 8'hfe; g = 8'hc3; b = 8'h95; end
	10'h228: begin r = 8'hfc; g = 8'hbb; b = 8'h85; end
	10'h248: begin r = 8'hf5; g = 8'hb8; b = 8'h7b; end
	10'h268: begin r = 8'hfb; g = 8'hbb; b = 8'h82; end
	10'h288: begin r = 8'hfd; g = 8'hc2; b = 8'h90; end
	10'h2a8: begin r = 8'hff; g = 8'hc3; b = 8'h98; end
	10'h2c8: begin r = 8'hfe; g = 8'hc9; b = 8'ha4; end
	10'h2e8: begin r = 8'hfe; g = 8'hce; b = 8'haa; end
	10'h308: begin r = 8'hec; g = 8'hba; b = 8'h8a; end
	10'h328: begin r = 8'hd8; g = 8'haa; b = 8'h74; end
	10'h348: begin r = 8'hc6; g = 8'hae; b = 8'h8e; end
	10'h368: begin r = 8'hae; g = 8'hb5; b = 8'haa; end
	10'h388: begin r = 8'h86; g = 8'ha9; b = 8'ha6; end
	10'h3a8: begin r = 8'h88; g = 8'ha6; b = 8'ha4; end
	10'h3c8: begin r = 8'h8d; g = 8'ha7; b = 8'ha6; end
	10'h3e8: begin r = 8'h89; g = 8'ha1; b = 8'ha1; end
	10'h009: begin r = 8'h9a; g = 8'hb4; b = 8'hb7; end
	10'h029: begin r = 8'h9b; g = 8'hb3; b = 8'hb3; end
	10'h049: begin r = 8'h9b; g = 8'hb4; b = 8'hb7; end
	10'h069: begin r = 8'h98; g = 8'hb5; b = 8'hb7; end
	10'h089: begin r = 8'h95; g = 8'hb3; b = 8'hb4; end
	10'h0a9: begin r = 8'h93; g = 8'h9d; b = 8'h98; end
	10'h0c9: begin r = 8'ha0; g = 8'h96; b = 8'h89; end
	10'h0e9: begin r = 8'ha0; g = 8'h85; b = 8'h5f; end
	10'h109: begin r = 8'hcc; g = 8'h97; b = 8'h3d; end
	10'h129: begin r = 8'hd1; g = 8'h9f; b = 8'h43; end
	10'h149: begin r = 8'hd3; g = 8'h9d; b = 8'h49; end
	10'h169: begin r = 8'hd9; g = 8'h9f; b = 8'h4d; end
	10'h189: begin r = 8'hdc; g = 8'ha4; b = 8'h52; end
	10'h1a9: begin r = 8'hdb; g = 8'ha5; b = 8'h5b; end
	10'h1c9: begin r = 8'hec; g = 8'hb6; b = 8'h79; end
	10'h1e9: begin r = 8'hfc; g = 8'hc6; b = 8'h99; end
	10'h209: begin r = 8'hf9; g = 8'hbe; b = 8'h8a; end
	10'h229: begin r = 8'hf0; g = 8'hb6; b = 8'h77; end
	10'h249: begin r = 8'hf0; g = 8'hb6; b = 8'h7a; end
	10'h269: begin r = 8'hf4; g = 8'hb8; b = 8'h7c; end
	10'h289: begin r = 8'hf7; g = 8'hba; b = 8'h82; end
	10'h2a9: begin r = 8'hf8; g = 8'hba; b = 8'h83; end
	10'h2c9: begin r = 8'hfd; g = 8'hc6; b = 8'h9a; end
	10'h2e9: begin r = 8'hff; g = 8'hd0; b = 8'hac; end
	10'h309: begin r = 8'hef; g = 8'hbb; b = 8'h8c; end
	10'h329: begin r = 8'hdc; g = 8'hac; b = 8'h7d; end
	10'h349: begin r = 8'hc8; g = 8'hac; b = 8'h84; end
	10'h369: begin r = 8'hb5; g = 8'hb4; b = 8'ha9; end
	10'h389: begin r = 8'h88; g = 8'haa; b = 8'ha8; end
	10'h3a9: begin r = 8'h87; g = 8'ha8; b = 8'ha5; end
	10'h3c9: begin r = 8'h89; g = 8'ha8; b = 8'ha6; end
	10'h3e9: begin r = 8'h88; g = 8'ha5; b = 8'ha3; end
	10'h00a: begin r = 8'h9c; g = 8'hb4; b = 8'hb7; end
	10'h02a: begin r = 8'h9c; g = 8'hb2; b = 8'hb3; end
	10'h04a: begin r = 8'h9c; g = 8'hb3; b = 8'hb5; end
	10'h06a: begin r = 8'h9a; g = 8'hb3; b = 8'hb5; end
	10'h08a: begin r = 8'h95; g = 8'hb3; b = 8'hb5; end
	10'h0aa: begin r = 8'h93; g = 8'ha1; b = 8'h95; end
	10'h0ca: begin r = 8'h8e; g = 8'h81; b = 8'h68; end
	10'h0ea: begin r = 8'ha7; g = 8'h8c; b = 8'h61; end
	10'h10a: begin r = 8'hc9; g = 8'h95; b = 8'h36; end
	10'h12a: begin r = 8'hce; g = 8'h99; b = 8'h3f; end
	10'h14a: begin r = 8'hd0; g = 8'h9a; b = 8'h45; end
	10'h16a: begin r = 8'hd7; g = 8'h9c; b = 8'h4b; end
	10'h18a: begin r = 8'hd6; g = 8'ha0; b = 8'h4d; end
	10'h1aa: begin r = 8'hda; g = 8'ha6; b = 8'h5b; end
	10'h1ca: begin r = 8'he4; g = 8'haf; b = 8'h6e; end
	10'h1ea: begin r = 8'hf1; g = 8'hb9; b = 8'h86; end
	10'h20a: begin r = 8'hee; g = 8'hb4; b = 8'h7d; end
	10'h22a: begin r = 8'he8; g = 8'hb1; b = 8'h6f; end
	10'h24a: begin r = 8'hed; g = 8'hb3; b = 8'h79; end
	10'h26a: begin r = 8'hea; g = 8'hb4; b = 8'h74; end
	10'h28a: begin r = 8'hec; g = 8'hb1; b = 8'h6c; end
	10'h2aa: begin r = 8'hee; g = 8'hb3; b = 8'h74; end
	10'h2ca: begin r = 8'hf1; g = 8'hb9; b = 8'h81; end
	10'h2ea: begin r = 8'hf0; g = 8'hbb; b = 8'h84; end
	10'h30a: begin r = 8'he3; g = 8'haf; b = 8'h74; end
	10'h32a: begin r = 8'hdd; g = 8'ha9; b = 8'h6e; end
	10'h34a: begin r = 8'hc8; g = 8'ha5; b = 8'h70; end
	10'h36a: begin r = 8'hb6; g = 8'hbb; b = 8'hae; end
	10'h38a: begin r = 8'h88; g = 8'hab; b = 8'ha7; end
	10'h3aa: begin r = 8'h85; g = 8'ha8; b = 8'ha4; end
	10'h3ca: begin r = 8'h88; g = 8'haa; b = 8'ha6; end
	10'h3ea: begin r = 8'h86; g = 8'ha7; b = 8'ha4; end
	10'h00b: begin r = 8'h9d; g = 8'hb5; b = 8'hb7; end
	10'h02b: begin r = 8'h9d; g = 8'hb3; b = 8'hb3; end
	10'h04b: begin r = 8'h9b; g = 8'hb1; b = 8'hb2; end
	10'h06b: begin r = 8'ha4; g = 8'hb2; b = 8'haa; end
	10'h08b: begin r = 8'hc8; g = 8'ha6; b = 8'h75; end
	10'h0ab: begin r = 8'ha4; g = 8'h98; b = 8'h81; end
	10'h0cb: begin r = 8'h8f; g = 8'h79; b = 8'h5f; end
	10'h0eb: begin r = 8'hb3; g = 8'h97; b = 8'h6d; end
	10'h10b: begin r = 8'hca; g = 8'h95; b = 8'h3a; end
	10'h12b: begin r = 8'hcd; g = 8'h9a; b = 8'h40; end
	10'h14b: begin r = 8'hcd; g = 8'h99; b = 8'h43; end
	10'h16b: begin r = 8'hd3; g = 8'h9b; b = 8'h45; end
	10'h18b: begin r = 8'hd4; g = 8'h9c; b = 8'h46; end
	10'h1ab: begin r = 8'hd9; g = 8'ha4; b = 8'h57; end
	10'h1cb: begin r = 8'heb; g = 8'hb2; b = 8'h75; end
	10'h1eb: begin r = 8'hf7; g = 8'hc0; b = 8'h98; end
	10'h20b: begin r = 8'hf4; g = 8'hbb; b = 8'h8d; end
	10'h22b: begin r = 8'hef; g = 8'hb8; b = 8'h80; end
	10'h24b: begin r = 8'he8; g = 8'hb3; b = 8'h76; end
	10'h26b: begin r = 8'he2; g = 8'hae; b = 8'h6d; end
	10'h28b: begin r = 8'he3; g = 8'haf; b = 8'h64; end
	10'h2ab: begin r = 8'he7; g = 8'hb0; b = 8'h6f; end
	10'h2cb: begin r = 8'hef; g = 8'hb8; b = 8'h7f; end
	10'h2eb: begin r = 8'hea; g = 8'hb6; b = 8'h7c; end
	10'h30b: begin r = 8'hdb; g = 8'ha8; b = 8'h64; end
	10'h32b: begin r = 8'hd9; g = 8'ha5; b = 8'h65; end
	10'h34b: begin r = 8'hc4; g = 8'ha1; b = 8'h6e; end
	10'h36b: begin r = 8'ha9; g = 8'hb0; b = 8'ha0; end
	10'h38b: begin r = 8'h85; g = 8'ha9; b = 8'ha6; end
	10'h3ab: begin r = 8'h86; g = 8'ha8; b = 8'ha9; end
	10'h3cb: begin r = 8'h85; g = 8'ha8; b = 8'ha5; end
	10'h3eb: begin r = 8'h83; g = 8'ha6; b = 8'ha2; end
	10'h00c: begin r = 8'h9e; g = 8'hb4; b = 8'hb6; end
	10'h02c: begin r = 8'h9f; g = 8'hb4; b = 8'hb6; end
	10'h04c: begin r = 8'h9d; g = 8'hb5; b = 8'hb8; end
	10'h06c: begin r = 8'hc8; g = 8'ha5; b = 8'h74; end
	10'h08c: begin r = 8'hd5; g = 8'h9e; b = 8'h53; end
	10'h0ac: begin r = 8'hcf; g = 8'ha2; b = 8'h5f; end
	10'h0cc: begin r = 8'ha9; g = 8'h98; b = 8'h79; end
	10'h0ec: begin r = 8'hb4; g = 8'h98; b = 8'h6b; end
	10'h10c: begin r = 8'hc9; g = 8'h9a; b = 8'h3d; end
	10'h12c: begin r = 8'hce; g = 8'h9d; b = 8'h48; end
	10'h14c: begin r = 8'hcd; g = 8'h98; b = 8'h42; end
	10'h16c: begin r = 8'hcb; g = 8'h94; b = 8'h39; end
	10'h18c: begin r = 8'hd0; g = 8'h99; b = 8'h3f; end
	10'h1ac: begin r = 8'hd9; g = 8'ha3; b = 8'h50; end
	10'h1cc: begin r = 8'hee; g = 8'hb4; b = 8'h79; end
	10'h1ec: begin r = 8'hf6; g = 8'hc1; b = 8'h8c; end
	10'h20c: begin r = 8'hfa; g = 8'hbc; b = 8'h88; end
	10'h22c: begin r = 8'hf8; g = 8'hbb; b = 8'h85; end
	10'h24c: begin r = 8'hf6; g = 8'hbe; b = 8'h85; end
	10'h26c: begin r = 8'hef; g = 8'hb7; b = 8'h79; end
	10'h28c: begin r = 8'hf1; g = 8'hb5; b = 8'h76; end
	10'h2ac: begin r = 8'hf3; g = 8'hb8; b = 8'h7c; end
	10'h2cc: begin r = 8'hf8; g = 8'hbc; b = 8'h81; end
	10'h2ec: begin r = 8'he8; g = 8'hb2; b = 8'h76; end
	10'h30c: begin r = 8'hd5; g = 8'ha2; b = 8'h57; end
	10'h32c: begin r = 8'hd6; g = 8'ha3; b = 8'h5a; end
	10'h34c: begin r = 8'hbc; g = 8'h9a; b = 8'h6a; end
	10'h36c: begin r = 8'h9d; g = 8'ha3; b = 8'h92; end
	10'h38c: begin r = 8'h82; g = 8'ha9; b = 8'ha5; end
	10'h3ac: begin r = 8'h82; g = 8'ha7; b = 8'ha7; end
	10'h3cc: begin r = 8'h83; g = 8'ha6; b = 8'ha2; end
	10'h3ec: begin r = 8'h82; g = 8'ha5; b = 8'ha1; end
	10'h00d: begin r = 8'h9e; g = 8'hb3; b = 8'hb7; end
	10'h02d: begin r = 8'h9d; g = 8'hb3; b = 8'hb6; end
	10'h04d: begin r = 8'h9c; g = 8'hb5; b = 8'hb6; end
	10'h06d: begin r = 8'hca; g = 8'h9d; b = 8'h5f; end
	10'h08d: begin r = 8'he7; g = 8'hae; b = 8'h6e; end
	10'h0ad: begin r = 8'hdc; g = 8'ha4; b = 8'h64; end
	10'h0cd: begin r = 8'hb1; g = 8'h9a; b = 8'h6b; end
	10'h0ed: begin r = 8'hb5; g = 8'h9d; b = 8'h70; end
	10'h10d: begin r = 8'hc7; g = 8'h98; b = 8'h49; end
	10'h12d: begin r = 8'hcf; g = 8'h9f; b = 8'h4d; end
	10'h14d: begin r = 8'hcc; g = 8'h98; b = 8'h3d; end
	10'h16d: begin r = 8'hca; g = 8'h94; b = 8'h39; end
	10'h18d: begin r = 8'hd1; g = 8'h99; b = 8'h41; end
	10'h1ad: begin r = 8'hdf; g = 8'haa; b = 8'h5f; end
	10'h1cd: begin r = 8'hf0; g = 8'hb7; b = 8'h7c; end
	10'h1ed: begin r = 8'hef; g = 8'hba; b = 8'h85; end
	10'h20d: begin r = 8'hf1; g = 8'hb7; b = 8'h77; end
	10'h22d: begin r = 8'hfb; g = 8'hbc; b = 8'h86; end
	10'h24d: begin r = 8'hf8; g = 8'hbe; b = 8'h86; end
	10'h26d: begin r = 8'hf7; g = 8'hb9; b = 8'h80; end
	10'h28d: begin r = 8'hf6; g = 8'hb8; b = 8'h7b; end
	10'h2ad: begin r = 8'hf9; g = 8'hba; b = 8'h82; end
	10'h2cd: begin r = 8'hf6; g = 8'hbc; b = 8'h83; end
	10'h2ed: begin r = 8'he9; g = 8'had; b = 8'h72; end
	10'h30d: begin r = 8'hd7; g = 8'ha3; b = 8'h58; end
	10'h32d: begin r = 8'hd1; g = 8'h9f; b = 8'h56; end
	10'h34d: begin r = 8'haf; g = 8'h92; b = 8'h61; end
	10'h36d: begin r = 8'h9a; g = 8'ha3; b = 8'h96; end
	10'h38d: begin r = 8'h81; g = 8'ha9; b = 8'ha5; end
	10'h3ad: begin r = 8'h81; g = 8'ha8; b = 8'ha7; end
	10'h3cd: begin r = 8'h83; g = 8'ha6; b = 8'ha2; end
	10'h3ed: begin r = 8'h81; g = 8'ha5; b = 8'ha1; end
	10'h00e: begin r = 8'h9c; g = 8'hb1; b = 8'hb4; end
	10'h02e: begin r = 8'h9d; g = 8'hb2; b = 8'hb5; end
	10'h04e: begin r = 8'h9b; g = 8'hb2; b = 8'hb6; end
	10'h06e: begin r = 8'hc9; g = 8'h9e; b = 8'h60; end
	10'h08e: begin r = 8'he8; g = 8'hac; b = 8'h63; end
	10'h0ae: begin r = 8'hb7; g = 8'h7d; b = 8'h1c; end
	10'h0ce: begin r = 8'hce; g = 8'h9f; b = 8'h56; end
	10'h0ee: begin r = 8'hb6; g = 8'h85; b = 8'h30; end
	10'h10e: begin r = 8'hcd; g = 8'h93; b = 8'h38; end
	10'h12e: begin r = 8'hd8; g = 8'ha0; b = 8'h4b; end
	10'h14e: begin r = 8'hd0; g = 8'h9b; b = 8'h42; end
	10'h16e: begin r = 8'hcb; g = 8'h98; b = 8'h44; end
	10'h18e: begin r = 8'hbe; g = 8'h8d; b = 8'h41; end
	10'h1ae: begin r = 8'haf; g = 8'h82; b = 8'h42; end
	10'h1ce: begin r = 8'h9d; g = 8'h6c; b = 8'h2a; end
	10'h1ee: begin r = 8'hc1; g = 8'h91; b = 8'h43; end
	10'h20e: begin r = 8'he6; g = 8'hb0; b = 8'h69; end
	10'h22e: begin r = 8'heb; g = 8'hb0; b = 8'h64; end
	10'h24e: begin r = 8'hef; g = 8'hb5; b = 8'h75; end
	10'h26e: begin r = 8'hec; g = 8'hb3; b = 8'h6c; end
	10'h28e: begin r = 8'hec; g = 8'hb0; b = 8'h6a; end
	10'h2ae: begin r = 8'hee; g = 8'hb3; b = 8'h76; end
	10'h2ce: begin r = 8'he8; g = 8'hae; b = 8'h6a; end
	10'h2ee: begin r = 8'hea; g = 8'hb1; b = 8'h6d; end
	10'h30e: begin r = 8'hdf; g = 8'haa; b = 8'h5c; end
	10'h32e: begin r = 8'hc8; g = 8'h99; b = 8'h4d; end
	10'h34e: begin r = 8'ha5; g = 8'h90; b = 8'h6f; end
	10'h36e: begin r = 8'h94; g = 8'ha5; b = 8'h99; end
	10'h38e: begin r = 8'h85; g = 8'ha9; b = 8'ha6; end
	10'h3ae: begin r = 8'h86; g = 8'ha8; b = 8'ha9; end
	10'h3ce: begin r = 8'h85; g = 8'ha7; b = 8'ha7; end
	10'h3ee: begin r = 8'h84; g = 8'ha7; b = 8'ha3; end
	10'h00f: begin r = 8'h9c; g = 8'hb2; b = 8'hb3; end
	10'h02f: begin r = 8'h9c; g = 8'hb1; b = 8'hb6; end
	10'h04f: begin r = 8'h9a; g = 8'hb0; b = 8'hb3; end
	10'h06f: begin r = 8'hb7; g = 8'ha6; b = 8'h82; end
	10'h08f: begin r = 8'hdc; g = 8'ha1; b = 8'h60; end
	10'h0af: begin r = 8'he3; g = 8'haa; b = 8'h67; end
	10'h0cf: begin r = 8'hc9; g = 8'h95; b = 8'h4a; end
	10'h0ef: begin r = 8'hbe; g = 8'h86; b = 8'h31; end
	10'h10f: begin r = 8'hd4; g = 8'h96; b = 8'h32; end
	10'h12f: begin r = 8'hdb; g = 8'ha1; b = 8'h3f; end
	10'h14f: begin r = 8'hdb; g = 8'ha2; b = 8'h4b; end
	10'h16f: begin r = 8'hd2; g = 8'h9e; b = 8'h55; end
	10'h18f: begin r = 8'hb3; g = 8'h84; b = 8'h3b; end
	10'h1af: begin r = 8'h8b; g = 8'h5d; b = 8'h20; end
	10'h1cf: begin r = 8'h81; g = 8'h58; b = 8'h26; end
	10'h1ef: begin r = 8'h8d; g = 8'h61; b = 8'h37; end
	10'h20f: begin r = 8'h9c; g = 8'h6a; b = 8'h19; end
	10'h22f: begin r = 8'hc5; g = 8'h8d; b = 8'h33; end
	10'h24f: begin r = 8'hd6; g = 8'ha2; b = 8'h4f; end
	10'h26f: begin r = 8'hd6; g = 8'ha2; b = 8'h55; end
	10'h28f: begin r = 8'hce; g = 8'h9b; b = 8'h4d; end
	10'h2af: begin r = 8'hd0; g = 8'h9e; b = 8'h53; end
	10'h2cf: begin r = 8'hd4; g = 8'ha4; b = 8'h65; end
	10'h2ef: begin r = 8'he0; g = 8'hae; b = 8'h72; end
	10'h30f: begin r = 8'hdb; g = 8'ha6; b = 8'h5a; end
	10'h32f: begin r = 8'hc4; g = 8'h92; b = 8'h42; end
	10'h34f: begin r = 8'hb5; g = 8'h9a; b = 8'h6c; end
	10'h36f: begin r = 8'h87; g = 8'haa; b = 8'ha5; end
	10'h38f: begin r = 8'h81; g = 8'ha9; b = 8'ha6; end
	10'h3af: begin r = 8'h86; g = 8'ha8; b = 8'ha8; end
	10'h3cf: begin r = 8'h85; g = 8'ha8; b = 8'ha4; end
	10'h3ef: begin r = 8'h84; g = 8'ha7; b = 8'ha3; end
	10'h010: begin r = 8'h9a; g = 8'hb2; b = 8'hb5; end
	10'h030: begin r = 8'h9c; g = 8'hb0; b = 8'hb4; end
	10'h050: begin r = 8'h9a; g = 8'hb0; b = 8'hb3; end
	10'h070: begin r = 8'ha5; g = 8'ha9; b = 8'ha1; end
	10'h090: begin r = 8'hdf; g = 8'ha2; b = 8'h59; end
	10'h0b0: begin r = 8'hdd; g = 8'ha3; b = 8'h59; end
	10'h0d0: begin r = 8'hd8; g = 8'h9f; b = 8'h56; end
	10'h0f0: begin r = 8'hbf; g = 8'h83; b = 8'h23; end
	10'h110: begin r = 8'hd1; g = 8'h92; b = 8'h27; end
	10'h130: begin r = 8'he5; g = 8'ha4; b = 8'h45; end
	10'h150: begin r = 8'hef; g = 8'hae; b = 8'h5e; end
	10'h170: begin r = 8'he7; g = 8'hab; b = 8'h60; end
	10'h190: begin r = 8'hd6; g = 8'ha0; b = 8'h59; end
	10'h1b0: begin r = 8'hcf; g = 8'ha4; b = 8'h75; end
	10'h1d0: begin r = 8'h90; g = 8'h72; b = 8'h41; end
	10'h1f0: begin r = 8'h86; g = 8'h63; b = 8'h39; end
	10'h210: begin r = 8'h75; g = 8'h50; b = 8'h1f; end
	10'h230: begin r = 8'hb3; g = 8'h83; b = 8'h30; end
	10'h250: begin r = 8'hd3; g = 8'ha1; b = 8'h52; end
	10'h270: begin r = 8'hb8; g = 8'h88; b = 8'h38; end
	10'h290: begin r = 8'h85; g = 8'h54; b = 8'h11; end
	10'h2b0: begin r = 8'h74; g = 8'h4e; b = 8'h1c; end
	10'h2d0: begin r = 8'h8c; g = 8'h64; b = 8'h2e; end
	10'h2f0: begin r = 8'ha2; g = 8'h77; b = 8'h39; end
	10'h310: begin r = 8'hba; g = 8'h8a; b = 8'h40; end
	10'h330: begin r = 8'hc6; g = 8'h90; b = 8'h42; end
	10'h350: begin r = 8'hb4; g = 8'h9b; b = 8'h64; end
	10'h370: begin r = 8'h88; g = 8'hab; b = 8'ha9; end
	10'h390: begin r = 8'h84; g = 8'haa; b = 8'ha6; end
	10'h3b0: begin r = 8'h85; g = 8'ha8; b = 8'ha4; end
	10'h3d0: begin r = 8'h85; g = 8'ha8; b = 8'ha4; end
	10'h3f0: begin r = 8'h84; g = 8'ha7; b = 8'ha3; end
	10'h011: begin r = 8'h9c; g = 8'hb1; b = 8'hb6; end
	10'h031: begin r = 8'h9b; g = 8'haf; b = 8'hb5; end
	10'h051: begin r = 8'h9a; g = 8'hb0; b = 8'hb0; end
	10'h071: begin r = 8'h9d; g = 8'haf; b = 8'had; end
	10'h091: begin r = 8'heb; g = 8'hac; b = 8'h6a; end
	10'h0b1: begin r = 8'he8; g = 8'hab; b = 8'h61; end
	10'h0d1: begin r = 8'hd4; g = 8'h9a; b = 8'h42; end
	10'h0f1: begin r = 8'hc2; g = 8'h82; b = 8'h1d; end
	10'h111: begin r = 8'hcd; g = 8'h8d; b = 8'h2a; end
	10'h131: begin r = 8'he4; g = 8'ha3; b = 8'h44; end
	10'h151: begin r = 8'hf6; g = 8'hb2; b = 8'h64; end
	10'h171: begin r = 8'hfd; g = 8'hbb; b = 8'h7f; end
	10'h191: begin r = 8'hef; g = 8'hb2; b = 8'h74; end
	10'h1b1: begin r = 8'he1; g = 8'ha9; b = 8'h5b; end
	10'h1d1: begin r = 8'hc7; g = 8'h93; b = 8'h36; end
	10'h1f1: begin r = 8'hb4; g = 8'h7d; b = 8'h29; end
	10'h211: begin r = 8'hd2; g = 8'h9f; b = 8'h5b; end
	10'h231: begin r = 8'he0; g = 8'ha5; b = 8'h5b; end
	10'h251: begin r = 8'hec; g = 8'hb4; b = 8'h74; end
	10'h271: begin r = 8'h9c; g = 8'h73; b = 8'h3f; end
	10'h291: begin r = 8'h5f; g = 8'h3e; b = 8'h19; end
	10'h2b1: begin r = 8'h60; g = 8'h46; b = 8'h22; end
	10'h2d1: begin r = 8'h5d; g = 8'h48; b = 8'h28; end
	10'h2f1: begin r = 8'h88; g = 8'h63; b = 8'h34; end
	10'h311: begin r = 8'hcb; g = 8'h93; b = 8'h45; end
	10'h331: begin r = 8'hca; g = 8'h93; b = 8'h3e; end
	10'h351: begin r = 8'ha6; g = 8'haa; b = 8'h8a; end
	10'h371: begin r = 8'h83; g = 8'hab; b = 8'ha6; end
	10'h391: begin r = 8'h82; g = 8'ha9; b = 8'ha4; end
	10'h3b1: begin r = 8'h83; g = 8'ha9; b = 8'ha4; end
	10'h3d1: begin r = 8'h85; g = 8'ha8; b = 8'ha4; end
	10'h3f1: begin r = 8'h83; g = 8'ha6; b = 8'ha2; end
	10'h012: begin r = 8'h9b; g = 8'haf; b = 8'hb4; end
	10'h032: begin r = 8'h9a; g = 8'haf; b = 8'hb4; end
	10'h052: begin r = 8'h9a; g = 8'hae; b = 8'hb0; end
	10'h072: begin r = 8'h99; g = 8'haf; b = 8'haf; end
	10'h092: begin r = 8'hd9; g = 8'ha7; b = 8'h61; end
	10'h0b2: begin r = 8'hf8; g = 8'hb4; b = 8'h69; end
	10'h0d2: begin r = 8'hd3; g = 8'h96; b = 8'h41; end
	10'h0f2: begin r = 8'hc5; g = 8'h83; b = 8'h21; end
	10'h112: begin r = 8'hcb; g = 8'h8b; b = 8'h29; end
	10'h132: begin r = 8'hde; g = 8'h9c; b = 8'h3f; end
	10'h152: begin r = 8'hf3; g = 8'haf; b = 8'h5c; end
	10'h172: begin r = 8'hfd; g = 8'hba; b = 8'h7c; end
	10'h192: begin r = 8'hfe; g = 8'hbd; b = 8'h83; end
	10'h1b2: begin r = 8'hf8; g = 8'hb7; b = 8'h75; end
	10'h1d2: begin r = 8'hf4; g = 8'hb2; b = 8'h6a; end
	10'h1f2: begin r = 8'hf6; g = 8'hb5; b = 8'h6b; end
	10'h212: begin r = 8'hf5; g = 8'hb2; b = 8'h6b; end
	10'h232: begin r = 8'he7; g = 8'ha5; b = 8'h50; end
	10'h252: begin r = 8'hf9; g = 8'hbb; b = 8'h87; end
	10'h272: begin r = 8'hef; g = 8'hb7; b = 8'h7e; end
	10'h292: begin r = 8'hd3; g = 8'ha1; b = 8'h6f; end
	10'h2b2: begin r = 8'hd3; g = 8'h9f; b = 8'h56; end
	10'h2d2: begin r = 8'he5; g = 8'hae; b = 8'h6b; end
	10'h2f2: begin r = 8'he6; g = 8'hac; b = 8'h64; end
	10'h312: begin r = 8'he9; g = 8'hae; b = 8'h68; end
	10'h332: begin r = 8'hca; g = 8'h9a; b = 8'h4c; end
	10'h352: begin r = 8'h8a; g = 8'hac; b = 8'ha7; end
	10'h372: begin r = 8'h87; g = 8'hab; b = 8'ha7; end
	10'h392: begin r = 8'h88; g = 8'hac; b = 8'ha8; end
	10'h3b2: begin r = 8'h82; g = 8'ha9; b = 8'ha4; end
	10'h3d2: begin r = 8'h83; g = 8'ha8; b = 8'ha4; end
	10'h3f2: begin r = 8'h83; g = 8'ha6; b = 8'ha2; end
	10'h013: begin r = 8'h9b; g = 8'hb0; b = 8'hb5; end
	10'h033: begin r = 8'h98; g = 8'had; b = 8'haf; end
	10'h053: begin r = 8'h99; g = 8'hac; b = 8'had; end
	10'h073: begin r = 8'h9a; g = 8'hac; b = 8'had; end
	10'h093: begin r = 8'hab; g = 8'ha8; b = 8'h9b; end
	10'h0b3: begin r = 8'hc9; g = 8'ha4; b = 8'h77; end
	10'h0d3: begin r = 8'hb7; g = 8'h91; b = 8'h4c; end
	10'h0f3: begin r = 8'hc3; g = 8'h86; b = 8'h23; end
	10'h113: begin r = 8'hc4; g = 8'h84; b = 8'h17; end
	10'h133: begin r = 8'hd4; g = 8'h94; b = 8'h2d; end
	10'h153: begin r = 8'he8; g = 8'ha5; b = 8'h4f; end
	10'h173: begin r = 8'hfc; g = 8'hb8; b = 8'h7b; end
	10'h193: begin r = 8'hfe; g = 8'hbd; b = 8'h7e; end
	10'h1b3: begin r = 8'hfc; g = 8'hb9; b = 8'h7a; end
	10'h1d3: begin r = 8'hf6; g = 8'hb5; b = 8'h75; end
	10'h1f3: begin r = 8'hf4; g = 8'hb2; b = 8'h6a; end
	10'h213: begin r = 8'hf2; g = 8'hb1; b = 8'h5f; end
	10'h233: begin r = 8'he5; g = 8'ha6; b = 8'h4c; end
	10'h253: begin r = 8'hf8; g = 8'hc1; b = 8'h8d; end
	10'h273: begin r = 8'hf6; g = 8'hbc; b = 8'h84; end
	10'h293: begin r = 8'hff; g = 8'hc7; b = 8'h9e; end
	10'h2b3: begin r = 8'hf4; g = 8'hbd; b = 8'h8d; end
	10'h2d3: begin r = 8'hf7; g = 8'hbf; b = 8'h8f; end
	10'h2f3: begin r = 8'hf6; g = 8'hbc; b = 8'h8c; end
	10'h313: begin r = 8'he7; g = 8'hab; b = 8'h65; end
	10'h333: begin r = 8'hc7; g = 8'ha0; b = 8'h64; end
	10'h353: begin r = 8'h86; g = 8'had; b = 8'ha9; end
	10'h373: begin r = 8'h86; g = 8'had; b = 8'ha8; end
	10'h393: begin r = 8'h87; g = 8'haa; b = 8'ha6; end
	10'h3b3: begin r = 8'h82; g = 8'ha9; b = 8'ha4; end
	10'h3d3: begin r = 8'h84; g = 8'ha8; b = 8'ha4; end
	10'h3f3: begin r = 8'h87; g = 8'haa; b = 8'ha6; end
	10'h014: begin r = 8'h9a; g = 8'hae; b = 8'hb0; end
	10'h034: begin r = 8'h98; g = 8'hac; b = 8'had; end
	10'h054: begin r = 8'h97; g = 8'hab; b = 8'hac; end
	10'h074: begin r = 8'h98; g = 8'hab; b = 8'hab; end
	10'h094: begin r = 8'h9b; g = 8'haa; b = 8'ha8; end
	10'h0b4: begin r = 8'ha1; g = 8'ha9; b = 8'ha3; end
	10'h0d4: begin r = 8'hb2; g = 8'h9a; b = 8'h6b; end
	10'h0f4: begin r = 8'hc3; g = 8'h86; b = 8'h24; end
	10'h114: begin r = 8'hc1; g = 8'h82; b = 8'h18; end
	10'h134: begin r = 8'hca; g = 8'h8a; b = 8'h20; end
	10'h154: begin r = 8'hda; g = 8'h9a; b = 8'h3d; end
	10'h174: begin r = 8'hea; g = 8'ha8; b = 8'h5b; end
	10'h194: begin r = 8'hef; g = 8'hae; b = 8'h59; end
	10'h1b4: begin r = 8'hee; g = 8'hac; b = 8'h58; end
	10'h1d4: begin r = 8'he0; g = 8'h9f; b = 8'h37; end
	10'h1f4: begin r = 8'hd1; g = 8'h90; b = 8'h2c; end
	10'h214: begin r = 8'he1; g = 8'ha3; b = 8'h51; end
	10'h234: begin r = 8'he6; g = 8'ha6; b = 8'h55; end
	10'h254: begin r = 8'hfc; g = 8'hc3; b = 8'h90; end
	10'h274: begin r = 8'heb; g = 8'haf; b = 8'h68; end
	10'h294: begin r = 8'hf0; g = 8'hb5; b = 8'h7f; end
	10'h2b4: begin r = 8'hfe; g = 8'hc4; b = 8'h99; end
	10'h2d4: begin r = 8'hfe; g = 8'hca; b = 8'ha2; end
	10'h2f4: begin r = 8'hf8; g = 8'hb9; b = 8'h87; end
	10'h314: begin r = 8'hdb; g = 8'ha0; b = 8'h51; end
	10'h334: begin r = 8'hb7; g = 8'ha4; b = 8'h79; end
	10'h354: begin r = 8'h88; g = 8'haf; b = 8'had; end
	10'h374: begin r = 8'h89; g = 8'hb0; b = 8'hae; end
	10'h394: begin r = 8'h86; g = 8'had; b = 8'haa; end
	10'h3b4: begin r = 8'h84; g = 8'haa; b = 8'ha5; end
	10'h3d4: begin r = 8'h86; g = 8'ha9; b = 8'ha6; end
	10'h3f4: begin r = 8'h87; g = 8'hab; b = 8'ha6; end
	10'h015: begin r = 8'h9a; g = 8'hae; b = 8'haf; end
	10'h035: begin r = 8'h99; g = 8'hac; b = 8'hac; end
	10'h055: begin r = 8'h99; g = 8'hab; b = 8'hac; end
	10'h075: begin r = 8'h98; g = 8'haa; b = 8'hab; end
	10'h095: begin r = 8'h99; g = 8'ha9; b = 8'haa; end
	10'h0b5: begin r = 8'ha8; g = 8'hb0; b = 8'ha7; end
	10'h0d5: begin r = 8'hb8; g = 8'h9b; b = 8'h6b; end
	10'h0f5: begin r = 8'hbc; g = 8'h85; b = 8'h1c; end
	10'h115: begin r = 8'hc7; g = 8'h8f; b = 8'h2c; end
	10'h135: begin r = 8'hbe; g = 8'h86; b = 8'h24; end
	10'h155: begin r = 8'hca; g = 8'h8e; b = 8'h25; end
	10'h175: begin r = 8'hd7; g = 8'h9a; b = 8'h33; end
	10'h195: begin r = 8'hd7; g = 8'h99; b = 8'h37; end
	10'h1b5: begin r = 8'hd0; g = 8'h90; b = 8'h28; end
	10'h1d5: begin r = 8'hbf; g = 8'h7f; b = 8'h20; end
	10'h1f5: begin r = 8'hd4; g = 8'h97; b = 8'h31; end
	10'h215: begin r = 8'hed; g = 8'hae; b = 8'h64; end
	10'h235: begin r = 8'heb; g = 8'had; b = 8'h64; end
	10'h255: begin r = 8'hfe; g = 8'hd1; b = 8'ha7; end
	10'h275: begin r = 8'hed; g = 8'hb3; b = 8'h74; end
	10'h295: begin r = 8'hc0; g = 8'h8a; b = 8'h35; end
	10'h2b5: begin r = 8'he7; g = 8'ha8; b = 8'h5e; end
	10'h2d5: begin r = 8'hf4; g = 8'hb2; b = 8'h71; end
	10'h2f5: begin r = 8'he8; g = 8'ha8; b = 8'h5e; end
	10'h315: begin r = 8'hd0; g = 8'h9a; b = 8'h49; end
	10'h335: begin r = 8'h99; g = 8'hab; b = 8'ha6; end
	10'h355: begin r = 8'h8e; g = 8'hb0; b = 8'hb0; end
	10'h375: begin r = 8'h8d; g = 8'haf; b = 8'hb0; end
	10'h395: begin r = 8'h8b; g = 8'haf; b = 8'haf; end
	10'h3b5: begin r = 8'h88; g = 8'hae; b = 8'hab; end
	10'h3d5: begin r = 8'h88; g = 8'hab; b = 8'ha7; end
	10'h3f5: begin r = 8'h88; g = 8'haa; b = 8'hab; end
	10'h016: begin r = 8'h9b; g = 8'had; b = 8'hae; end
	10'h036: begin r = 8'h98; g = 8'haa; b = 8'haa; end
	10'h056: begin r = 8'h98; g = 8'ha9; b = 8'ha9; end
	10'h076: begin r = 8'h99; g = 8'haa; b = 8'hab; end
	10'h096: begin r = 8'h9a; g = 8'haa; b = 8'ha7; end
	10'h0b6: begin r = 8'hbc; g = 8'hb4; b = 8'ha5; end
	10'h0d6: begin r = 8'hb3; g = 8'h9a; b = 8'h6a; end
	10'h0f6: begin r = 8'hba; g = 8'h83; b = 8'h28; end
	10'h116: begin r = 8'hc9; g = 8'h94; b = 8'h3b; end
	10'h136: begin r = 8'hb8; g = 8'h88; b = 8'h18; end
	10'h156: begin r = 8'hcc; g = 8'h91; b = 8'h35; end
	10'h176: begin r = 8'hcd; g = 8'h94; b = 8'h38; end
	10'h196: begin r = 8'hc0; g = 8'h85; b = 8'h29; end
	10'h1b6: begin r = 8'hb8; g = 8'h77; b = 8'h2a; end
	10'h1d6: begin r = 8'he9; g = 8'hac; b = 8'h6b; end
	10'h1f6: begin r = 8'hef; g = 8'hb0; b = 8'h6f; end
	10'h216: begin r = 8'hc7; g = 8'h89; b = 8'h33; end
	10'h236: begin r = 8'hdb; g = 8'h9c; b = 8'h4c; end
	10'h256: begin r = 8'he0; g = 8'ha9; b = 8'h60; end
	10'h276: begin r = 8'hd4; g = 8'ha1; b = 8'h5f; end
	10'h296: begin r = 8'h9b; g = 8'h5f; b = 8'h22; end
	10'h2b6: begin r = 8'hbe; g = 8'h7f; b = 8'h23; end
	10'h2d6: begin r = 8'hd3; g = 8'h95; b = 8'h2c; end
	10'h2f6: begin r = 8'hd3; g = 8'h92; b = 8'h28; end
	10'h316: begin r = 8'hca; g = 8'ha6; b = 8'h73; end
	10'h336: begin r = 8'hab; g = 8'hb1; b = 8'ha9; end
	10'h356: begin r = 8'h9f; g = 8'hb6; b = 8'hb4; end
	10'h376: begin r = 8'h91; g = 8'hb1; b = 8'hb0; end
	10'h396: begin r = 8'h8d; g = 8'hb2; b = 8'hb0; end
	10'h3b6: begin r = 8'h8b; g = 8'haf; b = 8'had; end
	10'h3d6: begin r = 8'h85; g = 8'had; b = 8'ha9; end
	10'h3f6: begin r = 8'h84; g = 8'ha9; b = 8'ha7; end
	10'h017: begin r = 8'h99; g = 8'haa; b = 8'hab; end
	10'h037: begin r = 8'h99; g = 8'ha9; b = 8'ha9; end
	10'h057: begin r = 8'h99; g = 8'ha8; b = 8'ha9; end
	10'h077: begin r = 8'h9b; g = 8'haa; b = 8'haa; end
	10'h097: begin r = 8'hab; g = 8'haf; b = 8'ha5; end
	10'h0b7: begin r = 8'hcf; g = 8'hc3; b = 8'haf; end
	10'h0d7: begin r = 8'h9b; g = 8'h76; b = 8'h4a; end
	10'h0f7: begin r = 8'hae; g = 8'h76; b = 8'h1b; end
	10'h117: begin r = 8'hc2; g = 8'h8e; b = 8'h2e; end
	10'h137: begin r = 8'hc0; g = 8'h8e; b = 8'h2c; end
	10'h157: begin r = 8'hcd; g = 8'h97; b = 8'h41; end
	10'h177: begin r = 8'hcf; g = 8'h9b; b = 8'h40; end
	10'h197: begin r = 8'hc0; g = 8'h87; b = 8'h3a; end
	10'h1b7: begin r = 8'he0; g = 8'ha7; b = 8'h55; end
	10'h1d7: begin r = 8'he5; g = 8'haa; b = 8'h5e; end
	10'h1f7: begin r = 8'hec; g = 8'hb0; b = 8'h6a; end
	10'h217: begin r = 8'he6; g = 8'haa; b = 8'h60; end
	10'h237: begin r = 8'hc2; g = 8'h89; b = 8'h2d; end
	10'h257: begin r = 8'hb0; g = 8'h79; b = 8'h24; end
	10'h277: begin r = 8'hcf; g = 8'h9e; b = 8'h55; end
	10'h297: begin r = 8'hb9; g = 8'h8f; b = 8'h4e; end
	10'h2b7: begin r = 8'ha8; g = 8'h6d; b = 8'h1f; end
	10'h2d7: begin r = 8'hcb; g = 8'h8f; b = 8'h24; end
	10'h2f7: begin r = 8'hd6; g = 8'ha0; b = 8'h48; end
	10'h317: begin r = 8'he2; g = 8'hc4; b = 8'h9f; end
	10'h337: begin r = 8'hda; g = 8'hcb; b = 8'hb5; end
	10'h357: begin r = 8'hd8; g = 8'hd1; b = 8'hc5; end
	10'h377: begin r = 8'hd5; g = 8'hd4; b = 8'hc7; end
	10'h397: begin r = 8'hc8; g = 8'hcf; b = 8'hc5; end
	10'h3b7: begin r = 8'hae; g = 8'hc1; b = 8'hbc; end
	10'h3d7: begin r = 8'h95; g = 8'hb1; b = 8'hb0; end
	10'h3f7: begin r = 8'h86; g = 8'hac; b = 8'ha6; end
	10'h018: begin r = 8'h9a; g = 8'ha9; b = 8'ha9; end
	10'h038: begin r = 8'h9a; g = 8'ha7; b = 8'ha6; end
	10'h058: begin r = 8'h9c; g = 8'ha8; b = 8'ha5; end
	10'h078: begin r = 8'h9f; g = 8'ha8; b = 8'h9d; end
	10'h098: begin r = 8'hce; g = 8'hc1; b = 8'had; end
	10'h0b8: begin r = 8'he8; g = 8'hda; b = 8'hc5; end
	10'h0d8: begin r = 8'h92; g = 8'h75; b = 8'h4a; end
	10'h0f8: begin r = 8'hbd; g = 8'h8a; b = 8'h2d; end
	10'h118: begin r = 8'hb4; g = 8'h7e; b = 8'h25; end
	10'h138: begin r = 8'hc2; g = 8'h90; b = 8'h37; end
	10'h158: begin r = 8'hce; g = 8'h98; b = 8'h41; end
	10'h178: begin r = 8'hd6; g = 8'ha3; b = 8'h50; end
	10'h198: begin r = 8'hd1; g = 8'h9d; b = 8'h49; end
	10'h1b8: begin r = 8'hc4; g = 8'h8b; b = 8'h2f; end
	10'h1d8: begin r = 8'hcb; g = 8'h93; b = 8'h44; end
	10'h1f8: begin r = 8'hcb; g = 8'h93; b = 8'h3e; end
	10'h218: begin r = 8'hd8; g = 8'h9c; b = 8'h43; end
	10'h238: begin r = 8'hd5; g = 8'ha0; b = 8'h4f; end
	10'h258: begin r = 8'hc3; g = 8'h92; b = 8'h3e; end
	10'h278: begin r = 8'hc4; g = 8'h95; b = 8'h36; end
	10'h298: begin r = 8'hba; g = 8'h89; b = 8'h41; end
	10'h2b8: begin r = 8'hb3; g = 8'h7e; b = 8'h31; end
	10'h2d8: begin r = 8'hda; g = 8'ha2; b = 8'h4b; end
	10'h2f8: begin r = 8'hd9; g = 8'hae; b = 8'h71; end
	10'h318: begin r = 8'hf3; g = 8'hdd; b = 8'hbc; end
	10'h338: begin r = 8'hd9; g = 8'hc9; b = 8'hb7; end
	10'h358: begin r = 8'hdf; g = 8'hd1; b = 8'hc1; end
	10'h378: begin r = 8'he3; g = 8'hd2; b = 8'hc4; end
	10'h398: begin r = 8'he3; g = 8'hd6; b = 8'hc7; end
	10'h3b8: begin r = 8'he2; g = 8'hdb; b = 8'hcb; end
	10'h3d8: begin r = 8'he1; g = 8'hdf; b = 8'hd1; end
	10'h3f8: begin r = 8'hb4; g = 8'hc2; b = 8'hba; end
	10'h019: begin r = 8'ha5; g = 8'had; b = 8'ha7; end
	10'h039: begin r = 8'hbd; g = 8'hbc; b = 8'hb0; end
	10'h059: begin r = 8'hcf; g = 8'hcb; b = 8'hbb; end
	10'h079: begin r = 8'hca; g = 8'hb9; b = 8'h99; end
	10'h099: begin r = 8'hdf; g = 8'hcc; b = 8'hbd; end
	10'h0b9: begin r = 8'he6; g = 8'hd6; b = 8'hc3; end
	10'h0d9: begin r = 8'he1; g = 8'hd2; b = 8'hb5; end
	10'h0f9: begin r = 8'hc0; g = 8'h87; b = 8'h2b; end
	10'h119: begin r = 8'hb4; g = 8'h80; b = 8'h28; end
	10'h139: begin r = 8'hb8; g = 8'h85; b = 8'h2c; end
	10'h159: begin r = 8'hc7; g = 8'h93; b = 8'h3c; end
	10'h179: begin r = 8'hce; g = 8'h9d; b = 8'h46; end
	10'h199: begin r = 8'hd4; g = 8'h9f; b = 8'h47; end
	10'h1b9: begin r = 8'hd2; g = 8'h9c; b = 8'h41; end
	10'h1d9: begin r = 8'he0; g = 8'ha5; b = 8'h54; end
	10'h1f9: begin r = 8'he7; g = 8'ha8; b = 8'h5f; end
	10'h219: begin r = 8'hde; g = 8'h9a; b = 8'h53; end
	10'h239: begin r = 8'hd8; g = 8'h97; b = 8'h47; end
	10'h259: begin r = 8'hd8; g = 8'h9a; b = 8'h49; end
	10'h279: begin r = 8'hdd; g = 8'ha1; b = 8'h50; end
	10'h299: begin r = 8'hd2; g = 8'ha0; b = 8'h54; end
	10'h2b9: begin r = 8'hca; g = 8'h95; b = 8'h49; end
	10'h2d9: begin r = 8'hd2; g = 8'h9e; b = 8'h4a; end
	10'h2f9: begin r = 8'he6; g = 8'hc4; b = 8'h9f; end
	10'h319: begin r = 8'hfb; g = 8'he2; b = 8'hc6; end
	10'h339: begin r = 8'hdb; g = 8'hcc; b = 8'hba; end
	10'h359: begin r = 8'hea; g = 8'hdb; b = 8'hc8; end
	10'h379: begin r = 8'hd5; g = 8'hc7; b = 8'hb5; end
	10'h399: begin r = 8'hdd; g = 8'hcf; b = 8'hbf; end
	10'h3b9: begin r = 8'hdb; g = 8'hcf; b = 8'hbf; end
	10'h3d9: begin r = 8'hf2; g = 8'he6; b = 8'hd4; end
	10'h3f9: begin r = 8'hdc; g = 8'hd2; b = 8'hc3; end
	10'h01a: begin r = 8'he0; g = 8'hd4; b = 8'hc0; end
	10'h03a: begin r = 8'hec; g = 8'he0; b = 8'hc7; end
	10'h05a: begin r = 8'hf4; g = 8'he6; b = 8'hcd; end
	10'h07a: begin r = 8'hdb; g = 8'hc8; b = 8'ha5; end
	10'h09a: begin r = 8'he1; g = 8'hd0; b = 8'hbc; end
	10'h0ba: begin r = 8'he3; g = 8'hd1; b = 8'hbf; end
	10'h0da: begin r = 8'hee; g = 8'hdd; b = 8'hc4; end
	10'h0fa: begin r = 8'he5; g = 8'hd0; b = 8'hab; end
	10'h11a: begin r = 8'hc2; g = 8'h91; b = 8'h3f; end
	10'h13a: begin r = 8'hae; g = 8'h7d; b = 8'h20; end
	10'h15a: begin r = 8'hbe; g = 8'h8e; b = 8'h3b; end
	10'h17a: begin r = 8'hc8; g = 8'h94; b = 8'h3f; end
	10'h19a: begin r = 8'hd1; g = 8'h9b; b = 8'h41; end
	10'h1ba: begin r = 8'he5; g = 8'had; b = 8'h5a; end
	10'h1da: begin r = 8'he7; g = 8'hab; b = 8'h59; end
	10'h1fa: begin r = 8'he7; g = 8'hab; b = 8'h58; end
	10'h21a: begin r = 8'hd7; g = 8'h9c; b = 8'h3b; end
	10'h23a: begin r = 8'hd1; g = 8'h91; b = 8'h35; end
	10'h25a: begin r = 8'hce; g = 8'h94; b = 8'h36; end
	10'h27a: begin r = 8'hdb; g = 8'ha4; b = 8'h4c; end
	10'h29a: begin r = 8'hde; g = 8'ha5; b = 8'h5a; end
	10'h2ba: begin r = 8'hce; g = 8'h9a; b = 8'h47; end
	10'h2da: begin r = 8'hd4; g = 8'haa; b = 8'h70; end
	10'h2fa: begin r = 8'hf2; g = 8'hd3; b = 8'hb3; end
	10'h31a: begin r = 8'hf6; g = 8'hde; b = 8'hc1; end
	10'h33a: begin r = 8'hdf; g = 8'hcf; b = 8'hbd; end
	10'h35a: begin r = 8'hf3; g = 8'he3; b = 8'hcf; end
	10'h37a: begin r = 8'hc9; g = 8'hb8; b = 8'ha7; end
	10'h39a: begin r = 8'hd1; g = 8'hc2; b = 8'hb2; end
	10'h3ba: begin r = 8'hd8; g = 8'hcc; b = 8'hbb; end
	10'h3da: begin r = 8'hee; g = 8'he1; b = 8'hcc; end
	10'h3fa: begin r = 8'hd4; g = 8'hc8; b = 8'hb8; end
	10'h01b: begin r = 8'hf1; g = 8'he4; b = 8'hca; end
	10'h03b: begin r = 8'hf2; g = 8'he3; b = 8'hc9; end
	10'h05b: begin r = 8'hf9; g = 8'he7; b = 8'hce; end
	10'h07b: begin r = 8'he7; g = 8'hd5; b = 8'hb2; end
	10'h09b: begin r = 8'hef; g = 8'hde; b = 8'hc4; end
	10'h0bb: begin r = 8'he6; g = 8'hd6; b = 8'hc2; end
	10'h0db: begin r = 8'he8; g = 8'hd8; b = 8'hbe; end
	10'h0fb: begin r = 8'hed; g = 8'hdb; b = 8'hc3; end
	10'h11b: begin r = 8'hef; g = 8'he0; b = 8'hc3; end
	10'h13b: begin r = 8'hc6; g = 8'h9d; b = 8'h5f; end
	10'h15b: begin r = 8'hb5; g = 8'h89; b = 8'h3b; end
	10'h17b: begin r = 8'hc0; g = 8'h90; b = 8'h3b; end
	10'h19b: begin r = 8'hca; g = 8'h96; b = 8'h3e; end
	10'h1bb: begin r = 8'hda; g = 8'ha3; b = 8'h4b; end
	10'h1db: begin r = 8'he7; g = 8'haa; b = 8'h50; end
	10'h1fb: begin r = 8'hec; g = 8'hab; b = 8'h4f; end
	10'h21b: begin r = 8'he7; g = 8'ha8; b = 8'h4b; end
	10'h23b: begin r = 8'hde; g = 8'h9f; b = 8'h43; end
	10'h25b: begin r = 8'hda; g = 8'ha1; b = 8'h45; end
	10'h27b: begin r = 8'he3; g = 8'ha9; b = 8'h58; end
	10'h29b: begin r = 8'hdc; g = 8'ha5; b = 8'h52; end
	10'h2bb: begin r = 8'hce; g = 8'h9d; b = 8'h4d; end
	10'h2db: begin r = 8'hd9; g = 8'hc4; b = 8'ha9; end
	10'h2fb: begin r = 8'he1; g = 8'hc9; b = 8'ha1; end
	10'h31b: begin r = 8'hf0; g = 8'hdf; b = 8'hbf; end
	10'h33b: begin r = 8'heb; g = 8'hdc; b = 8'hc4; end
	10'h35b: begin r = 8'hf7; g = 8'he4; b = 8'hd0; end
	10'h37b: begin r = 8'hc5; g = 8'hb5; b = 8'ha1; end
	10'h39b: begin r = 8'hc4; g = 8'hb4; b = 8'ha1; end
	10'h3bb: begin r = 8'hd7; g = 8'hc8; b = 8'hb6; end
	10'h3db: begin r = 8'hef; g = 8'he3; b = 8'hcb; end
	10'h3fb: begin r = 8'hd6; g = 8'hc8; b = 8'hb6; end
	10'h01c: begin r = 8'hfd; g = 8'hf1; b = 8'hd4; end
	10'h03c: begin r = 8'hfd; g = 8'hf0; b = 8'hd3; end
	10'h05c: begin r = 8'hfe; g = 8'hf0; b = 8'hd1; end
	10'h07c: begin r = 8'hfe; g = 8'hf0; b = 8'hcf; end
	10'h09c: begin r = 8'hd1; g = 8'hbd; b = 8'h8e; end
	10'h0bc: begin r = 8'hf3; g = 8'he1; b = 8'hc6; end
	10'h0dc: begin r = 8'hee; g = 8'hdd; b = 8'hc5; end
	10'h0fc: begin r = 8'hf1; g = 8'hde; b = 8'hc6; end
	10'h11c: begin r = 8'hee; g = 8'hdc; b = 8'hc3; end
	10'h13c: begin r = 8'hf2; g = 8'he2; b = 8'hc9; end
	10'h15c: begin r = 8'he1; g = 8'hca; b = 8'ha1; end
	10'h17c: begin r = 8'hb7; g = 8'h91; b = 8'h53; end
	10'h19c: begin r = 8'hba; g = 8'h90; b = 8'h38; end
	10'h1bc: begin r = 8'hca; g = 8'h98; b = 8'h3c; end
	10'h1dc: begin r = 8'hd5; g = 8'h9e; b = 8'h3c; end
	10'h1fc: begin r = 8'he6; g = 8'ha5; b = 8'h46; end
	10'h21c: begin r = 8'hf2; g = 8'hae; b = 8'h58; end
	10'h23c: begin r = 8'hf9; g = 8'hb5; b = 8'h65; end
	10'h25c: begin r = 8'hf4; g = 8'hb2; b = 8'h6b; end
	10'h27c: begin r = 8'hde; g = 8'ha6; b = 8'h51; end
	10'h29c: begin r = 8'hd8; g = 8'ha5; b = 8'h59; end
	10'h2bc: begin r = 8'he8; g = 8'hca; b = 8'ha6; end
	10'h2dc: begin r = 8'he8; g = 8'hd5; b = 8'hb6; end
	10'h2fc: begin r = 8'hcd; g = 8'hb9; b = 8'h8f; end
	10'h31c: begin r = 8'hf6; g = 8'he3; b = 8'hc6; end
	10'h33c: begin r = 8'hf2; g = 8'he2; b = 8'hc9; end
	10'h35c: begin r = 8'hf8; g = 8'he6; b = 8'hcd; end
	10'h37c: begin r = 8'hcd; g = 8'hbd; b = 8'ha7; end
	10'h39c: begin r = 8'hbc; g = 8'had; b = 8'h9a; end
	10'h3bc: begin r = 8'hd7; g = 8'hc6; b = 8'hb5; end
	10'h3dc: begin r = 8'hf0; g = 8'he1; b = 8'hca; end
	10'h3fc: begin r = 8'hda; g = 8'hcd; b = 8'hba; end
	10'h01d: begin r = 8'hff; g = 8'hf8; b = 8'hd8; end
	10'h03d: begin r = 8'hff; g = 8'hf5; b = 8'hd3; end
	10'h05d: begin r = 8'hff; g = 8'hf4; b = 8'hd0; end
	10'h07d: begin r = 8'hff; g = 8'hf5; b = 8'hd2; end
	10'h09d: begin r = 8'hef; g = 8'he5; b = 8'hb9; end
	10'h0bd: begin r = 8'hf4; g = 8'he2; b = 8'hba; end
	10'h0dd: begin r = 8'hfa; g = 8'he7; b = 8'hc7; end
	10'h0fd: begin r = 8'hf9; g = 8'he6; b = 8'hc9; end
	10'h11d: begin r = 8'hf6; g = 8'he4; b = 8'hc7; end
	10'h13d: begin r = 8'hf4; g = 8'he3; b = 8'hc3; end
	10'h15d: begin r = 8'hf6; g = 8'he0; b = 8'hc1; end
	10'h17d: begin r = 8'hee; g = 8'hd8; b = 8'hb7; end
	10'h19d: begin r = 8'hb9; g = 8'h97; b = 8'h60; end
	10'h1bd: begin r = 8'hb2; g = 8'h8b; b = 8'h46; end
	10'h1dd: begin r = 8'hc5; g = 8'h97; b = 8'h44; end
	10'h1fd: begin r = 8'hcc; g = 8'h94; b = 8'h3b; end
	10'h21d: begin r = 8'hd1; g = 8'h98; b = 8'h3a; end
	10'h23d: begin r = 8'hd3; g = 8'h99; b = 8'h3d; end
	10'h25d: begin r = 8'hd3; g = 8'h99; b = 8'h37; end
	10'h27d: begin r = 8'he1; g = 8'hb5; b = 8'h73; end
	10'h29d: begin r = 8'hf9; g = 8'he5; b = 8'hc4; end
	10'h2bd: begin r = 8'he7; g = 8'hcf; b = 8'hb0; end
	10'h2dd: begin r = 8'hf5; g = 8'hde; b = 8'hc0; end
	10'h2fd: begin r = 8'hf5; g = 8'he1; b = 8'hba; end
	10'h31d: begin r = 8'hea; g = 8'hd7; b = 8'hb2; end
	10'h33d: begin r = 8'hf6; g = 8'he8; b = 8'hce; end
	10'h35d: begin r = 8'hf8; g = 8'he9; b = 8'hd2; end
	10'h37d: begin r = 8'hda; g = 8'hcb; b = 8'hb6; end
	10'h39d: begin r = 8'hbc; g = 8'had; b = 8'h9a; end
	10'h3bd: begin r = 8'hd7; g = 8'hc6; b = 8'hb3; end
	10'h3dd: begin r = 8'hef; g = 8'he1; b = 8'hcc; end
	10'h3fd: begin r = 8'heb; g = 8'he1; b = 8'hcd; end
	10'h01e: begin r = 8'hff; g = 8'hf8; b = 8'hd8; end
	10'h03e: begin r = 8'hff; g = 8'hf5; b = 8'hd0; end
	10'h05e: begin r = 8'hff; g = 8'hf5; b = 8'hcf; end
	10'h07e: begin r = 8'hff; g = 8'hf6; b = 8'hd0; end
	10'h09e: begin r = 8'hff; g = 8'hf9; b = 8'hd7; end
	10'h0be: begin r = 8'he0; g = 8'hd2; b = 8'ha4; end
	10'h0de: begin r = 8'hff; g = 8'hf3; b = 8'hce; end
	10'h0fe: begin r = 8'hff; g = 8'hf0; b = 8'hcd; end
	10'h11e: begin r = 8'hfe; g = 8'hec; b = 8'hcb; end
	10'h13e: begin r = 8'hfc; g = 8'hea; b = 8'hc9; end
	10'h15e: begin r = 8'hfd; g = 8'he8; b = 8'hca; end
	10'h17e: begin r = 8'hfc; g = 8'he8; b = 8'hca; end
	10'h19e: begin r = 8'he8; g = 8'hd5; b = 8'hb7; end
	10'h1be: begin r = 8'hc6; g = 8'hb5; b = 8'h9f; end
	10'h1de: begin r = 8'hbc; g = 8'had; b = 8'h8d; end
	10'h1fe: begin r = 8'hc5; g = 8'hac; b = 8'h7f; end
	10'h21e: begin r = 8'hcb; g = 8'hb0; b = 8'h81; end
	10'h23e: begin r = 8'hca; g = 8'hb0; b = 8'h82; end
	10'h25e: begin r = 8'he7; g = 8'hcc; b = 8'hab; end
	10'h27e: begin r = 8'hfa; g = 8'he5; b = 8'hc7; end
	10'h29e: begin r = 8'hed; g = 8'hd9; b = 8'hb7; end
	10'h2be: begin r = 8'he9; g = 8'hd4; b = 8'hb6; end
	10'h2de: begin r = 8'hfb; g = 8'he3; b = 8'hc4; end
	10'h2fe: begin r = 8'hff; g = 8'hef; b = 8'hcd; end
	10'h31e: begin r = 8'he3; g = 8'hcf; b = 8'ha3; end
	10'h33e: begin r = 8'hfa; g = 8'he9; b = 8'hcf; end
	10'h35e: begin r = 8'hf6; g = 8'he8; b = 8'hd0; end
	10'h37e: begin r = 8'he2; g = 8'hd4; b = 8'hbf; end
	10'h39e: begin r = 8'hc1; g = 8'hb0; b = 8'h9e; end
	10'h3be: begin r = 8'hd3; g = 8'hc6; b = 8'hb1; end
	10'h3de: begin r = 8'hfc; g = 8'hf4; b = 8'hde; end
	10'h3fe: begin r = 8'hfd; g = 8'hf9; b = 8'he4; end
	10'h01f: begin r = 8'hfe; g = 8'hf9; b = 8'hd5; end
	10'h03f: begin r = 8'hff; g = 8'hf7; b = 8'hd0; end
	10'h05f: begin r = 8'hfe; g = 8'hf5; b = 8'hce; end
	10'h07f: begin r = 8'hff; g = 8'hf7; b = 8'hd0; end
	10'h09f: begin r = 8'hfe; g = 8'hf7; b = 8'hd4; end
	10'h0bf: begin r = 8'hf6; g = 8'hee; b = 8'hc7; end
	10'h0df: begin r = 8'hf0; g = 8'he6; b = 8'hb4; end
	10'h0ff: begin r = 8'hfe; g = 8'hfa; b = 8'hdb; end
	10'h11f: begin r = 8'hfc; g = 8'hf5; b = 8'hd8; end
	10'h13f: begin r = 8'hfe; g = 8'hf2; b = 8'hd0; end
	10'h15f: begin r = 8'hfd; g = 8'hee; b = 8'hcd; end
	10'h17f: begin r = 8'hfe; g = 8'hea; b = 8'hc8; end
	10'h19f: begin r = 8'hfb; g = 8'he6; b = 8'hc5; end
	10'h1bf: begin r = 8'he6; g = 8'hd2; b = 8'hb3; end
	10'h1df: begin r = 8'hbe; g = 8'hb1; b = 8'h93; end
	10'h1ff: begin r = 8'hcb; g = 8'hbc; b = 8'ha1; end
	10'h21f: begin r = 8'hdc; g = 8'hd1; b = 8'hb1; end
	10'h23f: begin r = 8'hda; g = 8'hcc; b = 8'had; end
	10'h25f: begin r = 8'hf5; g = 8'he5; b = 8'hc8; end
	10'h27f: begin r = 8'hd4; g = 8'hc5; b = 8'ha3; end
	10'h29f: begin r = 8'hde; g = 8'hcb; b = 8'hac; end
	10'h2bf: begin r = 8'hef; g = 8'hdb; b = 8'hbd; end
	10'h2df: begin r = 8'hfc; g = 8'he6; b = 8'hc3; end
	10'h2ff: begin r = 8'hfd; g = 8'he9; b = 8'hc6; end
	10'h31f: begin r = 8'he3; g = 8'hcf; b = 8'ha4; end
	10'h33f: begin r = 8'hf8; g = 8'he8; b = 8'hcb; end
	10'h35f: begin r = 8'hf3; g = 8'he5; b = 8'hca; end
	10'h37f: begin r = 8'he8; g = 8'hd9; b = 8'hc4; end
	10'h39f: begin r = 8'hcf; g = 8'hbf; b = 8'had; end
	10'h3bf: begin r = 8'hf3; g = 8'hea; b = 8'hd7; end
	10'h3df: begin r = 8'hff; g = 8'hfe; b = 8'hf0; end
	10'h3ff: begin r = 8'hfa; g = 8'hf8; b = 8'he5; end
endcase
end
endmodule
